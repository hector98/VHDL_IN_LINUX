LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TestBench IS
END TestBench;

ARCHITECTURE NOT_SELECT OF TestBench IS
		SIGNAL A_TB: STD_LOGIC := '0';
		SIGNAL Q_TB : STD_LOGIC;

		COMPONENT COMP_NOT_WITH_SELECT_01092023
				PORT(
						A : IN STD_LOGIC;
						Q : OUT STD_LOGIC
				);
		END COMPONENT;

BEGIN
		UUT : COMP_NOT_WITH_SELECT_01092023
		PORT MAP(
				A => A_TB,
				Q => Q_TB
		);

		STIM_PROC : PROCESS
		BEGIN
				A_TB <= '0';
				WAIT FOR 10 NS;

				A_TB <= '1';
				WAIT FOR 10 NS;

				WAIT;

		END PROCESS;
END NOT_SELECT;

