LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COMP_AND_WITH_SELECT_25082023 IS
		PORT(
		A:IN STD_LOGIC;
		B:IN STD_LOGIC;
		Q:OUT STD_LOGIC
		);
END COMP_AND_WITH_SELECT_25082023;

ARCHITECTURE COMP_AND_WITH_SELECT_25082023 OF COMP_AND_WITH_SELECT_25082023 IS
SIGNAL C:STD_LOGIC_VECTOR(1 DOWNTO 0);
BEGIN
		C <= A&B;
		WITH C SELECT 
				Q <= '0' WHEN "00",
					 '0' WHEN "01",
					 '0' WHEN "10",
					 '1' WHEN "11",
					 '0' WHEN OTHERS;
				
				--WHEN "00" => 
					--	Q <= '0';
				--WHEN "01" =>
						--Q <= '0';
				--WHEN "10" =>
						--Q <= '0';
				--WHEN "11" => 
						--Q <= '1';

END COMP_AND_WITH_SELECT_25082023;
