LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COMP_AND_WHEN_ELSE_25082023 IS
		PORT (
		A:IN STD_LOGIC;
		B:IN STD_LOGIC;
		Q:OUT STD_LOGIC
		);
END COMP_AND_WHEN_ELSE_25082023;

ARCHITECTURE COMP_AND_WHEN_ELSE_25082023 OF COMP_AND_WHEN_ELSE_25082023 IS
		signal c: std_logic_vector(1 downto 0);
BEGIN
		c <= a & b;
		Q <= '0' WHEN c = "00" ELSE
			 '0' WHEN c = "01" ELSE
			 '0' WHEN c = "10" ELSE
			 '1' WHEN c = "11" ELSE
			 '0';

END COMP_AND_WHEN_ELSE_25082023;
