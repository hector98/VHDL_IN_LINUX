-- ************************************************************************************************
-- Development name: Hector Manuel Barrios Barrios                                   
-- Operating System: GNU/Linux
                                
-- Kernel version: 6.1.0-13-amd64
                                  
-- ghdl version: -- GHDL 2.0.0 (Debian 2.0.0+dfsg-6.2) [Dunoon edition]
--  Compiled with GNAT Version: 12.2.0
--  mcode code generator
-- Written by Tristan Gingold.
-- 
-- Copyright (C) 2003 - 2022 Tristan Gingold.
-- GHDL is free software, covered by the GNU General Public License.  There is NO
-- warranty; not even for MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.
                                                           
-- date create: mié 15 nov 2023 12:57:50 CST
                                         
-- ************************************************************************************************

library ieee;
use ieee.std_logic_1164.all;

entity test is
        
       port(
			clk: in std_logic;
			a: in std_logic_vector (1 downto 0)

       );

end test;

architecture test of test is
-- Aqui van las señales

-- Y los components
        
begin
--Apartir de aqui va el codigo de tu programa

end test;
